module alu_16v(cc, result, valA, valB, op, sub, lr, arlo);
    input [15:0]  valA, valB;
    input [2:0]   op;
    input         sub, lr, arlo;

    output [3:0]  cc;
    output [15:0] result;



endmodule