module ksa_16b_top(Out, X, Y):

endmodule