`timescale 1ns/100ps

module alu_16b_tb;



endmodule;